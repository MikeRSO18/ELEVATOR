 LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY RAM16 IS

PORT(add:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
mode:IN STD_LOGIC;
Qram:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END RAM16 ;
ARCHITECTURE BEH123 OF RAM16 IS
SIGNAL P:STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
with add select
P<=
"0000" WHEN "0000",
"0001" WHEN "0001",
"0010" WHEN "0010",
"0011" WHEN "0011",
"0100" WHEN "0100",
"0101" WHEN "0101",
"0110" WHEN "0110",
"0111" WHEN "0111",
"1000" WHEN "1000",
"1001" WHEN "1001",
"1010" WHEN "1010",
"1011" WHEN "1011",
"0000" WHEN OTHERS;

process(mode)
begin
if(mode='0') then
Qram<=P;
else
Qram<="0000";
end if;
end process;
END BEH123;