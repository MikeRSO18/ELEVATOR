LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY mux_4pares IS

PORT(fil1,col1,f2,c2,f3,c3:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
SEL:IN STD_LOGIC_VECTOR(1 DOWNTO 0);
DOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END mux_4pares ;


ARCHITECTURE BEH123 OF mux_4pares IS

BEGIN
with SEL select
DOUT<=

fil1&col1 WHEN "00",
f2&c2 WHEN "01",
f3&c3 WHEN "10",
"ZZZZZZZZZZZZZZZZ" WHEN OTHERS;


END BEH123;